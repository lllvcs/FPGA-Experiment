LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY trans IS
    PORT (
        input : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        output : OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END ENTITY trans;

ARCHITECTURE behav OF trans IS
BEGIN
    PROCESS (input) BEGIN
        CASE input(3 DOWNTO 0) IS
            WHEN "0000" => output<="00000011" ; -- 0
            WHEN "0001" => output<="10011111" ; -- 1
            WHEN "0010" => output<="00100101" ; -- 2
            WHEN "0011" => output<="00001101" ; -- 3
            WHEN "0100" => output<="10011001" ; -- 4
            WHEN "0101" => output<="01001001" ; -- 5
            WHEN "0110" => output<="01000001" ; -- 6
            WHEN "0111" => output<="00011111" ; -- 7
            WHEN "1000" => output<="00000001" ; -- 8
            WHEN "1001" => output<="00010001" ; -- 9 
            WHEN OTHERS => output<="11111111" ; -- NULL;
        END CASE;
    END PROCESS;
END ARCHITECTURE behav;
